`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:35:59 11/13/2016 
// Design Name: 
// Module Name:    ALU 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU(
     input signed[31:0] A,
     input signed[31:0] B,
	  input [4:0] msb,
	  input [4:0] lsb,
     output reg signed [31:0] Out,//혷�����
	  output Overflow,
	  input [3:0] OP
    );
	/*assign Out = OP==0 ? A+B : (
					OP==1 ? A-B	: (
					OP==2 ? A|B	: (
					OP==3 ? A&B	: (
					B<<16 ))))	
					;*/
	wire [32:0] AddOut;
	wire [32:0] SubOut;
	assign AddOut = {A[31],A} + {B[31],B};
	assign SubOut = {A[31],A} - {B[31],B};
	assign Overflow = (~(AddOut[32] == AddOut[31])&&(OP == 0)) || 
							(~(SubOut[32] == SubOut[31])&&(OP == 1));
	always @(*) begin
		if (OP == 0) Out = AddOut[31:0];
		if (OP == 1) Out = SubOut[31:0];
		if (OP == 2) Out = A|B;
		if (OP == 3) Out = A&B;
		if (OP == 4) Out = {B[15:0],{16{1'b0}}};//����д{16{0}}���ᱻ��Ϊ�Ǻü���0��
		if (OP == 5) Out = B<<A[4:0]; //logic left
		if (OP == 6) Out = B>>A[4:0]; //logic right
		if (OP == 7) Out = A<B ? 1:0;
		if (OP == 8) Out = {1'b0,A}<{1'b0,B} ? 1:0;
		if (OP == 9) Out = 	A[4:0] == 0? {{0{B[31]}},B[31:0]} :
									A[4:0] == 1? {{1{B[31]}},B[31:1]} :
									A[4:0] == 2? {{2{B[31]}},B[31:2]} :
									A[4:0] == 3? {{3{B[31]}},B[31:3]} :
									A[4:0] == 4? {{4{B[31]}},B[31:4]} :
									A[4:0] == 5? {{5{B[31]}},B[31:5]} :
									A[4:0] == 6? {{6{B[31]}},B[31:6]} :
									A[4:0] == 7? {{7{B[31]}},B[31:7]} :
									A[4:0] == 8? {{8{B[31]}},B[31:8]} :
									A[4:0] == 9? {{9{B[31]}},B[31:9]} :
									A[4:0] == 10? {{10{B[31]}},B[31:10]} :
									A[4:0] == 11? {{11{B[31]}},B[31:11]} :
									A[4:0] == 12? {{12{B[31]}},B[31:12]} :
									A[4:0] == 13? {{13{B[31]}},B[31:13]} :
									A[4:0] == 14? {{14{B[31]}},B[31:14]} :
									A[4:0] == 15? {{15{B[31]}},B[31:15]} :
									A[4:0] == 16? {{16{B[31]}},B[31:16]} :
									A[4:0] == 17? {{17{B[31]}},B[31:17]} :
									A[4:0] == 18? {{18{B[31]}},B[31:18]} :
									A[4:0] == 19? {{19{B[31]}},B[31:19]} :
									A[4:0] == 20? {{20{B[31]}},B[31:20]} :
									A[4:0] == 21? {{21{B[31]}},B[31:21]} :
									A[4:0] == 22? {{22{B[31]}},B[31:22]} :
									A[4:0] == 23? {{23{B[31]}},B[31:23]} :
									A[4:0] == 24? {{24{B[31]}},B[31:24]} :
									A[4:0] == 25? {{25{B[31]}},B[31:25]} :
									A[4:0] == 26? {{26{B[31]}},B[31:26]} :
									A[4:0] == 27? {{27{B[31]}},B[31:27]} :
									A[4:0] == 28? {{28{B[31]}},B[31:28]} :
									A[4:0] == 29? {{29{B[31]}},B[31:29]} :
									A[4:0] == 30? {{30{B[31]}},B[31:30]} :
									A[4:0] == 31? {{31{B[31]}},B[31:31]} :
									{{32{B[31]}}};
		if (OP == 10) Out = A^B;
		if (OP == 11) Out = ~(A|B);					 
		if (OP == 12) Out = ((B>>(msb+1) )<<(msb+1))|(( A<<(31-msb+lsb) )>>(31-msb))|((B << 32-lsb) >> (32-lsb));
		if (OP == 13) Out = (A << (31-msb-lsb)) >> (31-msb);
	end
endmodule
